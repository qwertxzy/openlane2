VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_256x16
  FOREIGN fakeram130_256x16 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 285.660 BY 187.680 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 5.850 0.800 6.150 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.250 0.800 8.550 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.650 0.800 10.950 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.050 0.800 13.350 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 15.450 0.800 15.750 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.850 0.800 18.150 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.250 0.800 20.550 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.650 0.800 22.950 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.050 0.800 25.350 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.450 0.800 27.750 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.850 0.800 30.150 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 32.250 0.800 32.550 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 34.650 0.800 34.950 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.050 0.800 37.350 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.450 0.800 39.750 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 41.850 0.800 42.150 ;
    END
  END w_mask_in[15]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 50.250 0.800 50.550 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.650 0.800 52.950 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.050 0.800 55.350 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 57.450 0.800 57.750 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.850 0.800 60.150 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 62.250 0.800 62.550 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 64.650 0.800 64.950 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.050 0.800 67.350 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 69.450 0.800 69.750 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.850 0.800 72.150 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.250 0.800 74.550 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.650 0.800 76.950 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 79.050 0.800 79.350 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.450 0.800 81.750 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 83.850 0.800 84.150 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 86.250 0.800 86.550 ;
    END
  END rd_out[15]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 94.650 0.800 94.950 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.050 0.800 97.350 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.450 0.800 99.750 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 101.850 0.800 102.150 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 104.250 0.800 104.550 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 106.650 0.800 106.950 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 109.050 0.800 109.350 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 111.450 0.800 111.750 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 113.850 0.800 114.150 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 116.250 0.800 116.550 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 118.650 0.800 118.950 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 121.050 0.800 121.350 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.450 0.800 123.750 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 125.850 0.800 126.150 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 128.250 0.800 128.550 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 130.650 0.800 130.950 ;
    END
  END wd_in[15]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.050 0.800 139.350 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 141.450 0.800 141.750 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 143.850 0.800 144.150 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 146.250 0.800 146.550 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.650 0.800 148.950 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 151.050 0.800 151.350 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 153.450 0.800 153.750 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 155.850 0.800 156.150 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 164.250 0.800 164.550 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 166.650 0.800 166.950 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.050 0.800 169.350 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 5.400 6.000 6.600 181.680 ;
      RECT 15.000 6.000 16.200 181.680 ;
      RECT 24.600 6.000 25.800 181.680 ;
      RECT 34.200 6.000 35.400 181.680 ;
      RECT 43.800 6.000 45.000 181.680 ;
      RECT 53.400 6.000 54.600 181.680 ;
      RECT 63.000 6.000 64.200 181.680 ;
      RECT 72.600 6.000 73.800 181.680 ;
      RECT 82.200 6.000 83.400 181.680 ;
      RECT 91.800 6.000 93.000 181.680 ;
      RECT 101.400 6.000 102.600 181.680 ;
      RECT 111.000 6.000 112.200 181.680 ;
      RECT 120.600 6.000 121.800 181.680 ;
      RECT 130.200 6.000 131.400 181.680 ;
      RECT 139.800 6.000 141.000 181.680 ;
      RECT 149.400 6.000 150.600 181.680 ;
      RECT 159.000 6.000 160.200 181.680 ;
      RECT 168.600 6.000 169.800 181.680 ;
      RECT 178.200 6.000 179.400 181.680 ;
      RECT 187.800 6.000 189.000 181.680 ;
      RECT 197.400 6.000 198.600 181.680 ;
      RECT 207.000 6.000 208.200 181.680 ;
      RECT 216.600 6.000 217.800 181.680 ;
      RECT 226.200 6.000 227.400 181.680 ;
      RECT 235.800 6.000 237.000 181.680 ;
      RECT 245.400 6.000 246.600 181.680 ;
      RECT 255.000 6.000 256.200 181.680 ;
      RECT 264.600 6.000 265.800 181.680 ;
      RECT 274.200 6.000 275.400 181.680 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 10.200 6.000 11.400 181.680 ;
      RECT 19.800 6.000 21.000 181.680 ;
      RECT 29.400 6.000 30.600 181.680 ;
      RECT 39.000 6.000 40.200 181.680 ;
      RECT 48.600 6.000 49.800 181.680 ;
      RECT 58.200 6.000 59.400 181.680 ;
      RECT 67.800 6.000 69.000 181.680 ;
      RECT 77.400 6.000 78.600 181.680 ;
      RECT 87.000 6.000 88.200 181.680 ;
      RECT 96.600 6.000 97.800 181.680 ;
      RECT 106.200 6.000 107.400 181.680 ;
      RECT 115.800 6.000 117.000 181.680 ;
      RECT 125.400 6.000 126.600 181.680 ;
      RECT 135.000 6.000 136.200 181.680 ;
      RECT 144.600 6.000 145.800 181.680 ;
      RECT 154.200 6.000 155.400 181.680 ;
      RECT 163.800 6.000 165.000 181.680 ;
      RECT 173.400 6.000 174.600 181.680 ;
      RECT 183.000 6.000 184.200 181.680 ;
      RECT 192.600 6.000 193.800 181.680 ;
      RECT 202.200 6.000 203.400 181.680 ;
      RECT 211.800 6.000 213.000 181.680 ;
      RECT 221.400 6.000 222.600 181.680 ;
      RECT 231.000 6.000 232.200 181.680 ;
      RECT 240.600 6.000 241.800 181.680 ;
      RECT 250.200 6.000 251.400 181.680 ;
      RECT 259.800 6.000 261.000 181.680 ;
      RECT 269.400 6.000 270.600 181.680 ;
      RECT 279.000 6.000 280.200 181.680 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 285.660 187.680 ;
    LAYER met2 ;
    RECT 0 0 285.660 187.680 ;
    LAYER met3 ;
    RECT 0.800 0 285.660 187.680 ;
    RECT 0 0.000 0.800 5.850 ;
    RECT 0 6.150 0.800 8.250 ;
    RECT 0 8.550 0.800 10.650 ;
    RECT 0 10.950 0.800 13.050 ;
    RECT 0 13.350 0.800 15.450 ;
    RECT 0 15.750 0.800 17.850 ;
    RECT 0 18.150 0.800 20.250 ;
    RECT 0 20.550 0.800 22.650 ;
    RECT 0 22.950 0.800 25.050 ;
    RECT 0 25.350 0.800 27.450 ;
    RECT 0 27.750 0.800 29.850 ;
    RECT 0 30.150 0.800 32.250 ;
    RECT 0 32.550 0.800 34.650 ;
    RECT 0 34.950 0.800 37.050 ;
    RECT 0 37.350 0.800 39.450 ;
    RECT 0 39.750 0.800 41.850 ;
    RECT 0 42.150 0.800 50.250 ;
    RECT 0 50.550 0.800 52.650 ;
    RECT 0 52.950 0.800 55.050 ;
    RECT 0 55.350 0.800 57.450 ;
    RECT 0 57.750 0.800 59.850 ;
    RECT 0 60.150 0.800 62.250 ;
    RECT 0 62.550 0.800 64.650 ;
    RECT 0 64.950 0.800 67.050 ;
    RECT 0 67.350 0.800 69.450 ;
    RECT 0 69.750 0.800 71.850 ;
    RECT 0 72.150 0.800 74.250 ;
    RECT 0 74.550 0.800 76.650 ;
    RECT 0 76.950 0.800 79.050 ;
    RECT 0 79.350 0.800 81.450 ;
    RECT 0 81.750 0.800 83.850 ;
    RECT 0 84.150 0.800 86.250 ;
    RECT 0 86.550 0.800 94.650 ;
    RECT 0 94.950 0.800 97.050 ;
    RECT 0 97.350 0.800 99.450 ;
    RECT 0 99.750 0.800 101.850 ;
    RECT 0 102.150 0.800 104.250 ;
    RECT 0 104.550 0.800 106.650 ;
    RECT 0 106.950 0.800 109.050 ;
    RECT 0 109.350 0.800 111.450 ;
    RECT 0 111.750 0.800 113.850 ;
    RECT 0 114.150 0.800 116.250 ;
    RECT 0 116.550 0.800 118.650 ;
    RECT 0 118.950 0.800 121.050 ;
    RECT 0 121.350 0.800 123.450 ;
    RECT 0 123.750 0.800 125.850 ;
    RECT 0 126.150 0.800 128.250 ;
    RECT 0 128.550 0.800 130.650 ;
    RECT 0 130.950 0.800 139.050 ;
    RECT 0 139.350 0.800 141.450 ;
    RECT 0 141.750 0.800 143.850 ;
    RECT 0 144.150 0.800 146.250 ;
    RECT 0 146.550 0.800 148.650 ;
    RECT 0 148.950 0.800 151.050 ;
    RECT 0 151.350 0.800 153.450 ;
    RECT 0 153.750 0.800 155.850 ;
    RECT 0 156.150 0.800 164.250 ;
    RECT 0 164.550 0.800 166.650 ;
    RECT 0 166.950 0.800 169.050 ;
    RECT 0 169.350 0.800 187.680 ;
    LAYER met4 ;
    RECT 0 0 285.660 6.000 ;
    RECT 0 181.680 285.660 187.680 ;
    RECT 0.000 6.000 5.400 181.680 ;
    RECT 6.600 6.000 10.200 181.680 ;
    RECT 11.400 6.000 15.000 181.680 ;
    RECT 16.200 6.000 19.800 181.680 ;
    RECT 21.000 6.000 24.600 181.680 ;
    RECT 25.800 6.000 29.400 181.680 ;
    RECT 30.600 6.000 34.200 181.680 ;
    RECT 35.400 6.000 39.000 181.680 ;
    RECT 40.200 6.000 43.800 181.680 ;
    RECT 45.000 6.000 48.600 181.680 ;
    RECT 49.800 6.000 53.400 181.680 ;
    RECT 54.600 6.000 58.200 181.680 ;
    RECT 59.400 6.000 63.000 181.680 ;
    RECT 64.200 6.000 67.800 181.680 ;
    RECT 69.000 6.000 72.600 181.680 ;
    RECT 73.800 6.000 77.400 181.680 ;
    RECT 78.600 6.000 82.200 181.680 ;
    RECT 83.400 6.000 87.000 181.680 ;
    RECT 88.200 6.000 91.800 181.680 ;
    RECT 93.000 6.000 96.600 181.680 ;
    RECT 97.800 6.000 101.400 181.680 ;
    RECT 102.600 6.000 106.200 181.680 ;
    RECT 107.400 6.000 111.000 181.680 ;
    RECT 112.200 6.000 115.800 181.680 ;
    RECT 117.000 6.000 120.600 181.680 ;
    RECT 121.800 6.000 125.400 181.680 ;
    RECT 126.600 6.000 130.200 181.680 ;
    RECT 131.400 6.000 135.000 181.680 ;
    RECT 136.200 6.000 139.800 181.680 ;
    RECT 141.000 6.000 144.600 181.680 ;
    RECT 145.800 6.000 149.400 181.680 ;
    RECT 150.600 6.000 154.200 181.680 ;
    RECT 155.400 6.000 159.000 181.680 ;
    RECT 160.200 6.000 163.800 181.680 ;
    RECT 165.000 6.000 168.600 181.680 ;
    RECT 169.800 6.000 173.400 181.680 ;
    RECT 174.600 6.000 178.200 181.680 ;
    RECT 179.400 6.000 183.000 181.680 ;
    RECT 184.200 6.000 187.800 181.680 ;
    RECT 189.000 6.000 192.600 181.680 ;
    RECT 193.800 6.000 197.400 181.680 ;
    RECT 198.600 6.000 202.200 181.680 ;
    RECT 203.400 6.000 207.000 181.680 ;
    RECT 208.200 6.000 211.800 181.680 ;
    RECT 213.000 6.000 216.600 181.680 ;
    RECT 217.800 6.000 221.400 181.680 ;
    RECT 222.600 6.000 226.200 181.680 ;
    RECT 227.400 6.000 231.000 181.680 ;
    RECT 232.200 6.000 235.800 181.680 ;
    RECT 237.000 6.000 240.600 181.680 ;
    RECT 241.800 6.000 245.400 181.680 ;
    RECT 246.600 6.000 250.200 181.680 ;
    RECT 251.400 6.000 255.000 181.680 ;
    RECT 256.200 6.000 259.800 181.680 ;
    RECT 261.000 6.000 264.600 181.680 ;
    RECT 265.800 6.000 269.400 181.680 ;
    RECT 270.600 6.000 274.200 181.680 ;
    RECT 275.400 6.000 279.000 181.680 ;
    RECT 280.200 6.000 285.660 181.680 ;
    LAYER OVERLAP ;
    RECT 0 0 285.660 187.680 ;
  END
END fakeram130_256x16

END LIBRARY
